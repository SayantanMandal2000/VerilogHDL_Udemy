module inverter(x,y);
  input x;
  output y;
  assign y=~x;
endmodule
